* C:\Users\Administrator\Documents\circuit\Schematic6.sch

* Schematics Version 9.1 - Web Update 1
* Thu Sep 02 19:30:27 2021



** Analysis setup **
.tran 0ns 1000ns
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic6.net"
.INC "Schematic6.als"


.probe


.END
